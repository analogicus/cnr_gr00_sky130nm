*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNRG00_IFT_lpe.spi
#else
.include ../../../work/xsch/CNRG00_IFT.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  0 dc {AVDD}

VPWR PWRUP_1V8 0 dc {AVDD}

.nodeset v(VDA) = 0.9
.nodeset v(VD) = 0.9
.nodeset v(LPI) = 0.9

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDA IBP4 IBP3 IBP2 IBP1 IBP0 VDD_1V8 VSS PWRUP_1V8 VD LPI LPI CNRG00_IFT

VIB4 IBP4 0 dc 0.9
VIB3 IBP3 0 dc 0.9
VIB2 IBP2 0 dc 0.9
VIBP1 IBP1 0 dc 0.9
VIBP0 IBP0 0 dc 0.9

B5 temp 0 v=temper

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save v(VDA) v(VD) v(IBP) v(VDD_1V8) v(VSS) v(PWRUP_1V8)

.save i(VIBP2) i(VIBP1) i(VIBP0)
.save v(temp)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100n 20u 0

dc TEMP -40 125 10
write
quit

.endc

.end
