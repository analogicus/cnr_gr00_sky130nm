*CNRG00 LSTB
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNRG00_IFT_lpe.spi
#else
.include ../../../work/xsch/CNRG00_IFT.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option reltol=1e-5 gmin=1e-15


*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  0  dc {AVDD}
VPWR  PWRUP_1V8  VSS  dc {AVDD}

*-----------------------------------------------------------------
* Loop stability
*-----------------------------------------------------------------
.include ../../../../cpdk/ngspice/tian_subckt.lib
X999 LPI LPO loopgainprobe

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDA IBP4 IBP3 IBP2 IBP1 IBP0 VDD_1V8 VSS PWRUP_1V8 VD LPO LPI CNRG00_IFT

*-----------------------------------------------------------------
* STASH
*-----------------------------------------------------------------
V4 IBP4 0 dc {AVDD/2}
V3 IBP3 0 dc {AVDD/2}
V2 IBP2 0 dc {AVDD/2}
V1 IBP1 0 dc {AVDD/2}
V0 IBP0 0 dc {AVDD/2}

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save V(X999.x) I(v.X999.Vi)
.save v(LPO) v(LPI) v(vd) v(vda)

#ifdef Debug
*.save all
#else


#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100n 20u 0
op
write {cicname}_op.raw

*----------------------------------------------------------------
* LSTB analysis
*----------------------------------------------------------------
* Set voltage AC to 1
ac dec 50 100 10G

* Set Current to 1
alter i.X999.Ii acmag=1
alter v.X999.Vi acmag=0
ac dec 50 100 10G

let lg_mag = db(tian_loop())
let lg_phase = 180*cph(tian_loop())/pi

*set gnuplot_terminal=png/quit
*gnuplot {cicname}_loop_gain lg_mag
*gnuplot {cicname}_loop_phase lg_phase

write

#ifdef Debug
*quit
#else

quit
#endif
.endc
