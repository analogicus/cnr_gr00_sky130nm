*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_GR00_lpe.spi
#else
.include ../../../work/lpe/SUNTR_CAP_20_lpe.spi
.include ../../../work/xsch/CNR_GR00.spice

#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-4

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

*- 8 MHz clock frequency
.param PERIOD_CLK = 100n

*- 25% duty-cycle clock
.param PW_CLK = PERIOD_CLK/2

*- Frequency bin of the input signal
.param fbin = 5

*- number of cycles in FFT
.param nbpt = 128

*- Sampling frequency
.param fs = 1/PERIOD_CLK

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  0  pwl 0 0 10n {AVDD}
VPW  PWRUP_1V8 0  pwl 0 0 10n {AVDD}
VRE  RESET_1V8 0   pwl 0 {AVDD} 1u {AVDD} 1.001u 0
VDWN  DOWN_N_1V8 0   pwl 0 {AVDD} 2u {AVDD} 2.001u 0

VCLK CK_1V8 0 dc 0 pulse (0 {AVDD} 1u {TRF} {TRF} {PW_CLK} {PERIOD_CLK})

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD_1V8 VSS PWRUP_1V8 RESET_1V8 VO_1V8 DO_1V8 CK_1V8 DO_1V8 CNR_GR00

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save v(VDD_1V8) v(VSS) v(PWRUP_1V8) v(RESET_1V8) v(VO_1V8) v(DOWN_N_1V8) v(DO_1V8) v(CK_1V8)
.save v(xdut.ibp) v(xdut.vd) v(xdut.vda) v(xdut.xt.vg) v(xdut.xt.voa) v(xdut.xt.vref)
.save v(xdut.xt.xota.vbp)
.save v(xdut.xt.xota.vbn1)
.save v(xdut.xt.xota.vbn2)
.save v(xdut.von) v(xdut.vop)
.save v(xdut.xcmp.von0)
.save v(xdut.xcmp.vop0)
.save v(xdut.xcmp.vs)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100p 2n 0

foreach vtemp -40 -20 0 20 40 80 125
  option temp=$vtemp
  tran 1n 20u 1n
  write {cicname}_$vtemp
end

quit


.endc

.end
