*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_GR00_lpe.spi
#else
.include ../../../work/lpe/SUNTR_CAP_20_lpe.spi
.include ../../../work/xsch/CNR_GR00.spice

#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-4

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 100p

.param t_start = 4u
.param t_start_del = {t_start + TRF}

*- 8 MHz clock frequency
.param PERIOD_CLK = 200n

*- 25% duty-cycle clock
.param PW_CLK = PERIOD_CLK/2

*- Supply, vdda is set in includes
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  0  dc {AVDD}
VPW  PWRUP_1V8 0  dc {AVDD}
VRE  RESET_1V8 0   pwl 0 {AVDD} {t_start} {AVDD} {t_start_del} 0

VCLK CK_1V8 0 dc 0 pulse 0 {AVDD} {t_start} {TRF} {TRF} {PW_CLK} {PERIOD_CLK}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD_1V8 VSS PWRUP_1V8 RESET_1V8 DO_1V8 CK_1V8 CNR_GR00

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save v(VDD_1V8) v(VSS) v(PWRUP_1V8) v(RESET_1V8)  v(DO_1V8) v(CK_1V8)
.save v(xdut.ibp) v(xdut.vd) v(xdut.vda) (xdut.vdb) v(xdut.xt.vg) v(xdut.xt.voa) v(xdut.xt.vref)
.save v(xdut.xt.xota.vbp)
.save v(xdut.xt.xota.vbn1)
.save v(xdut.xt.xota.vbn2)
.save v(xdut.vo)
.save v(xdut.vdb)
.save v(xdut.xi.vdb_on_1v8)
.save v(xdut.xi.vda_on_1v8)
.save v(xdut.xd.vop)
.save v(xdut.xd.von)
.save v(xdut.xd.xcmp.von0)
.save v(xdut.xd.xcmp.vop0)
.save v(xdut.xd.xcmp.vs)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100n 20u 0

#ifdef Nosweep


foreach vtemp -40 125
  option temp=$vtemp
  tran 1n 8u 1n
  write {cicname}_$vtemp
end

#else

foreach vtemp -40 -20 0 20 40 80 125
  option temp=$vtemp
*- 32*200n = 8.4 us =>
*- 64*200n = 16.8us => +5us =22us
  tran 1n 22u 1n
*- 128*200n = 25.6us => +5u = 31us
*- 256*200n = 55.2us => +5us = 61us
*  tran 1n 61u 1n
  write {cicname}_$vtemp
end

#endif

quit


.endc

.end
